/*
    This layer proceeds dense_0  
*/