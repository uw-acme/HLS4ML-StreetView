/*
    this layer proceeds bn_conv2d_2  
*/