/*
    This layer proceeds pooling_1  
*/