/*
    This is the initial conv2d layer after the input layer
*/