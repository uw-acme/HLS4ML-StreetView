/*
    This layer proceeds dense_1  
*/