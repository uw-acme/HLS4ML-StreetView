/*
    This layer proceeds dense_act_1 
*/ 