/*
    This layer proceeds bn_conv2d_1  
*/