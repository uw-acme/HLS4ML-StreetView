/*
    This layer proceeds bn_dense_0  
*/