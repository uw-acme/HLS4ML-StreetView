/*
    This layer proceeds flatten
*/