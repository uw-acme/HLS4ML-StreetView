/*
    this layer proceeds conv_act_1  
*/