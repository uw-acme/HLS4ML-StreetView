/*
    This layer proceeds conv2d_1  
*/