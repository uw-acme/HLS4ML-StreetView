/*
    This layer proceeds conv_act_2  
*/