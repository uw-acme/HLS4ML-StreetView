/*
    This layer proceeds ouput_dense  
*/