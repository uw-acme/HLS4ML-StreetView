/*
    this layer proceeds the pool_1
*/