/*
    This layer proceeds pool_2  
*/